grammar edu:umn:cs:melt:exts:ableC:unification:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:datatype:concretesyntax;
exports edu:umn:cs:melt:exts:ableC:algebraicDataTypes:patternmatching:concretesyntax;
exports edu:umn:cs:melt:exts:ableC:templating:concretesyntax;
exports edu:umn:cs:melt:exts:ableC:templateAlgebraicDataTypes:datatype:concretesyntax;
exports edu:umn:cs:melt:exts:ableC:string:concretesyntax;
exports edu:umn:cs:melt:exts:ableC:vector:concretesyntax;
exports edu:umn:cs:melt:exts:ableC:constructor:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:unification:concretesyntax:unification;
exports edu:umn:cs:melt:exts:ableC:unification:concretesyntax:allocation;
exports edu:umn:cs:melt:exts:ableC:unification:concretesyntax:patternmatching;
grammar edu:umn:cs:melt:exts:ableC:unification:concretesyntax:unification;

exports edu:umn:cs:melt:exts:ableC:string:concretesyntax;
